module top_module (
    input clk,
    input reset,
    input enable,
    output [3:0] Q,
    output c_enable,
    output c_load,
    output [3:0] c_d
); //
    assign c_enable = enable;
    always @(posedge clk) begin
        if (reset | Q == 12) begin
            c_load <= 0 ;
            c_d <= 1;  
        end
        else begin
            c_load <= 1;
        end
    end

    count4 the_counter (clk, c_enable, c_load, c_d, Q);

endmodule